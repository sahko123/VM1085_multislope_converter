-- spi_bus.vhd

-- Generated using ACDS version 22.1 915

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity spi_bus is
	port (
		ncs : in  std_logic := '0'; -- ncs.ncs
		osc : out std_logic;        -- osc.osc
		sck : in  std_logic := '0'; -- sck.sck
		si  : in  std_logic := '0'; --  si.si
		so  : out std_logic         --  so.so
	);
end entity spi_bus;

architecture rtl of spi_bus is
	component spi_bus_ufm_spi_0 is
		port (
			si  : in  std_logic := 'X'; -- si
			sck : in  std_logic := 'X'; -- sck
			ncs : in  std_logic := 'X'; -- ncs
			so  : out std_logic;        -- so
			osc : out std_logic         -- osc
		);
	end component spi_bus_ufm_spi_0;

begin

	ufm_spi_0 : component spi_bus_ufm_spi_0
		port map (
			si  => si,  --  si.si
			sck => sck, -- sck.sck
			ncs => ncs, -- ncs.ncs
			so  => so,  --  so.so
			osc => osc  -- osc.osc
		);

end architecture rtl; -- of spi_bus
