
module spi_bus (
	si,
	sck,
	ncs,
	so,
	osc);	

	input		si;
	input		sck;
	input		ncs;
	output		so;
	output		osc;
endmodule
