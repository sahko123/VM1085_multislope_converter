-- parallel_bus.vhd

-- Generated using ACDS version 22.1 915

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity parallel_bus is
	port (
		addr       : in  std_logic_vector(7 downto 0) := (others => '0'); --       addr.addr
		data_valid : out std_logic;                                       -- data_valid.data_valid
		datain     : in  std_logic_vector(7 downto 0) := (others => '0'); --     datain.datain
		dataout    : out std_logic_vector(7 downto 0);                    --    dataout.dataout
		nbusy      : out std_logic;                                       --      nbusy.nbusy
		nerase     : in  std_logic                    := '0';             --     nerase.nerase
		nread      : in  std_logic                    := '0';             --      nread.nread
		nwrite     : in  std_logic                    := '0';             --     nwrite.nwrite
		osc        : out std_logic                                        --        osc.osc
	);
end entity parallel_bus;

architecture rtl of parallel_bus is
	component parallel_bus_ufm_parallel_0 is
		port (
			addr       : in  std_logic_vector(7 downto 0) := (others => 'X'); -- addr
			nread      : in  std_logic                    := 'X';             -- nread
			dataout    : out std_logic_vector(7 downto 0);                    -- dataout
			nbusy      : out std_logic;                                       -- nbusy
			data_valid : out std_logic;                                       -- data_valid
			datain     : in  std_logic_vector(7 downto 0) := (others => 'X'); -- datain
			nwrite     : in  std_logic                    := 'X';             -- nwrite
			nerase     : in  std_logic                    := 'X';             -- nerase
			osc        : out std_logic                                        -- osc
		);
	end component parallel_bus_ufm_parallel_0;

begin

	ufm_parallel_0 : component parallel_bus_ufm_parallel_0
		port map (
			addr       => addr,       --       addr.addr
			nread      => nread,      --      nread.nread
			dataout    => dataout,    --    dataout.dataout
			nbusy      => nbusy,      --      nbusy.nbusy
			data_valid => data_valid, -- data_valid.data_valid
			datain     => datain,     --     datain.datain
			nwrite     => nwrite,     --     nwrite.nwrite
			nerase     => nerase,     --     nerase.nerase
			osc        => osc         --        osc.osc
		);

end architecture rtl; -- of parallel_bus
